library ieee;
use ieee.std_logic_1164.all;

----------------------------------------

entity Driver is
port(	x: in std_logic;
	F: out std_logic
);
end Driver;  

----------------------------------------
