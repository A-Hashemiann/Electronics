library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity Inverter is
    port (
        A : in  std_logic;  -- Input signal
        Y : out std_logic   -- Output signal
    );
end entity Inverter;